mstein19@remus.amherst.edu.49858:1471142699