mstein19@remus.amherst.edu.20072:1471142699