lschmidlein19@remus.amherst.edu.61859:1471142699