mstein19@remus.amherst.edu.49825:1471142699