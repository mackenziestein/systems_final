lschmidlein19@remus.amherst.edu.10533:1471142699